`ifndef ENVIRONMENT__SV
`define ENVIRONMENT__SV

`include "ethpack_generator.sv"
`include "driver2xgmii.sv"
`include "monitor4xgmii.sv"
`include "config.sv"
`include "scoreboard_pack.sv"

/////////////////////////////////////////////////////////
// Call scoreboard from Driver using callbacks
/////////////////////////////////////////////////////////
class Scb_Driver_cbs #(parameter XGMII_WIDTH = 64) extends Driver2xgmii_cbs #(.XGMII_WIDTH(XGMII_WIDTH));
    Scoreboard scb;

    function new(Scoreboard scb);
        this.scb = scb;
    endfunction

    // Send received pack to scoreboard
    virtual task post_tx(input Driver2xgmii #(.XGMII_WIDTH(XGMII_WIDTH)) drv, input Ethpack pack);
        scb.save_expected(pack);
    endtask
endclass 

/////////////////////////////////////////////////////////
// Call scoreboard from Monitor using callbacks
/////////////////////////////////////////////////////////
class Scb_Monitor_cbs #(parameter XGMII_WIDTH = 64) extends Monitor4xgmii_cbs #(.XGMII_WIDTH(XGMII_WIDTH));
    Scoreboard scb;

    function new(Scoreboard scb);
        this.scb = scb;
    endfunction

    // Send received cell to scoreboard
    virtual task post_rx(input Monitor4xgmii #(.XGMII_WIDTH(XGMII_WIDTH)) mon, input Ethpack pack);
        scb.check_actual(pack);
    endtask
endclass 

class Environment #(parameter XGMII_WIDTH_PMA = 32);
    Ethpack_generator genPma  [];
    mailbox genPma2drvPma     [];
    event   drvPma2genPma     [];
    Driver2xgmii  #(.XGMII_WIDTH(XGMII_WIDTH_PMA  )) drvPma  [];
    Monitor4xgmii #(.XGMII_WIDTH(XGMII_WIDTH_PMA  )) monPma  [];
    Config cfg;
    Scoreboard scb[];
    virtual xgmii_if#(XGMII_WIDTH_PMA  ).TbTx pmaTx;
    virtual xgmii_if#(XGMII_WIDTH_PMA  ).TbRx pmaRx;

    extern function new(input virtual xgmii_if#(XGMII_WIDTH_PMA  ).TbTx pmaTx, 
                        input virtual xgmii_if#(XGMII_WIDTH_PMA  ).TbRx pmaRx);
    extern virtual function void build();
    extern virtual task run();
    extern virtual task force_linkdown_pma();
    extern virtual function void wrap_up();

endclass

function Environment::new
    (
        input virtual xgmii_if#(XGMII_WIDTH_PMA  ).TbTx pmaTx,
        input virtual xgmii_if#(XGMII_WIDTH_PMA  ).TbRx pmaRx
    );

    this.pmaTx = pmaTx;
    this.pmaRx = pmaRx;

    cfg = new();
endfunction

function void Environment::build();

    genPma    = new[1];
    drvPma    = new[1];
    genPma2drvPma     = new[1];
    drvPma2genPma     = new[1];
    scb = new[1];
    scb[0] = new(cfg,"pma2pma");

    genPma2drvPma    [0] = new();
    genPma           [0] = new(genPma2drvPma    [0], drvPma2genPma    [0], cfg , "pma");
    drvPma           [0] = new(genPma2drvPma    [0], drvPma2genPma    [0], cfg,  pmaTx, 32, 1, "pma");

    monPma    = new[1];
    monPma   [0] = new(pmaRx, "pma");


    // Connect the scoreboard with callbacks
    begin
        Scb_Driver_cbs   #(.XGMII_WIDTH(XGMII_WIDTH_PMA  )) sdcPma    = new(scb[0]);
        Scb_Monitor_cbs  #(.XGMII_WIDTH(XGMII_WIDTH_PMA  )) smcPma    = new(scb[0]);
        foreach (drvPma  [i] ) drvPma[i].cbsq.push_back(sdcPma);  // Add scb to every driver
        foreach (monPma  [i] ) monPma[i].cbsq.push_back(smcPma);  // Add scb to every monitor
    end

endfunction

task Environment::run();
    
    int num_genPma_running;
    num_genPma_running = 1;

    foreach(genPma[i]) begin
        int j=i;      // Automatic variable to hold index in spawned threads
        fork begin
            genPma[j].run();       // Wait for generator to finish
            num_genPma_running--;  // Decrement driver count
        end
        drvPma[j].run();
        join_none
    end

    if (cfg.test_force_linkdown==1) begin
        fork begin
            this.force_linkdown_pma();
        end
        join_none
    end

    foreach(monPma[i]) begin
        int j=i;       // Automatic variable to hold index in spawned threads
        fork
            monPma[j].run();
        join_none
    end

    // Wait for all generators to finish, or time-out
    fork : timeout_block
        wait ((num_genPma_running == 0));
        begin
            repeat (1000000) @pmaTx.tbtx_cb;
            $display("@%0t: %m Env: ERROR: Timeout while waiting for generators to finish", $time);
            cfg.nErrors = cfg.nErrors + 1;
        end
    join_any
    disable timeout_block;

    // Wait a little longer for the data flow through switch, into monitors, and scoreboards
    repeat (1000) @pmaTx.tbtx_cb;

endtask : run

task Environment::force_linkdown_pma();
    int pause;
    int linkdown;
    forever begin
        @drvPma2genPma[0];
        pause = $urandom_range(500,600);
        linkdown = $urandom_range(200,300);
        repeat (pause) @pmaTx.tbtx_cb;
        top.dut_u.force_linkdown_pma = 1;
        repeat (linkdown) @pmaTx.tbtx_cb;
        top.dut_u.force_linkdown_pma = 0;
    end 
endtask

function void Environment::wrap_up();
    scb[0].wrap_up;
    $display("@%0t: Env: End of simulation, %0d ERROR, %0d WARNING", $time, cfg.nErrors, cfg.nWarnings);
endfunction

`endif 

